//####################################################################
//  Author: Austin | @SV-Engineer
//    Date: 28OCT2023
// Purpose: This header file is used to import all packages related
//          i2c RTL at once.
//####################################################################

`ifndef I2C_INCLUDE_SVH_
  `define I2C_INCLUDE_SVH_
  import i2c_primitives_pkg::*;
`endif /* I2C_INCLUDE_SVH_ */
