//####################################################################
//  Author: Austin | @SV-Engineer
//    Date: 29JUL2023
// Purpose: This file is for demonstrating threads and how we can use
//          events for adding some synchronicity.
//####################################################################

program unit_test (interface top_if);
  // This initial block will be the "main" thread that drives the rest.
  initial
    begin : main
    
    end : main


endprogram : unit_test
