//####################################################################
//  Author: Austin | @SV-Engineer
//    Date: 28OCT2023
// Purpose: This package is for defining some of the primitives
//          related to the i2c rtl.
//####################################################################

  // Section comment template
  // ========================
  // START - 
  // ========================

  // ========================
  // END - 
  // ========================

package i2c_primitives_pkg;

endpackage : i2c_primitives_pkg
