//####################################################################
//  Author: Austin | @SV-Engineer
//    Date: 28OCT2023
// Purpose: This header file is used to import all packages related
//          to the framework at once.
//####################################################################

`ifndef FRAME_WORK_SVH_
  `define FRAME_WORK_SVH_

  import primitives_pkg::*;

`endif /* FRAME_WORK_SVH_ */